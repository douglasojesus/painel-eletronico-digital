module Demultiplexador();

endmodule