library verilog;
use verilog.vl_types.all;
entity Letreiro_vlg_vec_tst is
end Letreiro_vlg_vec_tst;
