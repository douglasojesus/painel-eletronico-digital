module Letreiro(CLK, ch0, ch1, C1L1, C2L1, C3L1, C4L1, C5L1, C6L1, C7L1, C1L2, C2L2, C3L2, C4L2, C5L2, C6L2, C7L2, C1L3, C2L3, C3L3, C4L3, C5L3, C6L3, C7L3, C1L4, C2L4, C3L4, C4L4, C5L4, C6L4, C7L4, C1L5, C2L5, C3L5, C4L5, C5L5, C6L5, C7L5);

	input CLK, ch0, ch1;
	output C1L1, C2L1, C3L1, C4L1, C5L1, C6L1, C7L1;
	output C1L2, C2L2, C3L2, C4L2, C5L2, C6L2, C7L2;
	output C1L3, C2L3, C3L3, C4L3, C5L3, C6L3, C7L3;
	output C1L4, C2L4, C3L4, C4L4, C5L4, C6L4, C7L4;
	output C1L5, C2L5, C3L5, C4L5, C5L5, C6L5, C7L5;


		/*reg [15:0] L1 = 16'b1010_1110_1110_1110;
		reg [15:0] L2 = 16'b1010_1000_1000_1000;
		reg [15:0] L3 = 16'b1010_1110_1110_1110;
		reg [15:0] L4 = 16'b1010_1000_1000_0010;
		reg [15:0] L5 = 16'b1110_1110_1000_1110;*/
	
	RegistradorL1 instL1(ch0, ch1, CLK, C1L1, C2L1, C3L1, C4L1, C5L1, C6L1, C7L1);
	RegistradorL2 instL2(ch0, ch1, CLK, C1L2, C2L2, C3L2, C4L2, C5L2, C6L2, C7L2);
	RegistradorL3 instL3(ch0, ch1, CLK, C1L3, C2L3, C3L3, C4L3, C5L3, C6L3, C7L3);
  
endmodule
