library verilog;
use verilog.vl_types.all;
entity Letreiro_vlg_check_tst is
    port(
        C1              : in     vl_logic;
        C2              : in     vl_logic;
        C3              : in     vl_logic;
        C4              : in     vl_logic;
        C5              : in     vl_logic;
        C6              : in     vl_logic;
        C7              : in     vl_logic;
        L1              : in     vl_logic;
        L2              : in     vl_logic;
        L3              : in     vl_logic;
        L4              : in     vl_logic;
        L5              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Letreiro_vlg_check_tst;
